library verilog;
use verilog.vl_types.all;
entity MLP_FPGA_vlg_vec_tst is
end MLP_FPGA_vlg_vec_tst;
